<svg id="wave" style="transform:rotate(180deg)" 
viewBox="0 -5 1440 200" version="1.1" xmlns="http://www.w3.org/2000/svg"><defs>
<linearGradient id="sw-gradient-0" x1="0" x2="0" y1="0" y2="0">
<stop stop-color="rgba(254, 226, 213, 1)" offset="0%"></stop><stop stop-color="rgba(254, 226, 213, 1)" offset="100%"></stop>
</linearGradient></defs><path style="transform:translate(0, 0px); opacity:1" fill="url(#sw-gradient-0)" 
d="M0,20L40,26.7C80,33,160,47,240,60C320,73,400,87,480,106.7C560,127,640,153,720,146.7C800,140,880,100,960,83.3C1040,67,1120,73
,1200,83.3C1280,93,1360,107,1440,120C1520,133,1600,147,1680,130C1760,113,1840,67,1920,60C2000,53,2080,87,2160,106.7C2240,127,2320
,133,2400,116.7C2480,100,2560,60,2640,66.7C2720,73,2800,127,2880,133.3C2960,140,3040,100,3120,73.3C3200,47,3280,33,3360,40C3440
,47,3520,73,3600,73.3C3680,73,3760,47,3840,30C3920,13,4000,7,4080,33.3C4160,60,4240,120,4320,133.3C4400,147,4480,113,4560,106.7C4640,
100,4720,120,4800,116.7C4880,113,4960,87,5040,70C5120,53,5200,47,5280,40C5360,33,5440,27,5520,33.3C5600,40,5680,60,5720,70L5760,80L5760,
200L5720,200C5680,200,5600,200,5520,200C5440,200,5360,200,5280,200C5200,200,5120,200,5040,200C4960,200,4880,200,4800,200C4720,200,4640,
200,4560,200C4480,200,4400,200,4320,200C4240,200,4160,200,4080,200C4000,200,3920,200,3840,200C3760,200,3680,200,3600,200C3520,200,3440,
200,3360,200C3280,200,3200,200,3120,200C3040,200,2960,200,2880,200C2800,200,2720,200,2640,200C2560,200,2480,200,2400,200C2320,200,2240,
200,2160,200C2080,200,2000,200,1920,200C1840,200,1760,200,1680,200C1600,200,1520,200,1440,200C1360,200,1280,200,1200,200C1120,200,1040,
200,960,200C880,200,800,200,720,200C640,200,560,200,480,200C400,200,320,200,240,200C160,200,80,200,40,200L0,200Z"></path></svg>